* linguist-detectable
*.vhd linguist-language=VHDL
*.xml linguist-language=ignore
